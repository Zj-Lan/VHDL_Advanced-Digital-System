----------------------------------------------------------------------------------
-- Company: 	Artesis
-- Engineer: 	Kaj Van der Hallen
-- 
-- Create Date:    00:27:27 04/18/2012 
-- Module Name:    prom_DMH - Behavioral 
-- Project Name: Multifunctionele klok
-- Target Devices: FPGA
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity prom_DMH is
    Port ( clk : in std_logic;
			  addr : in std_logic_vector(8 downto 0);
           M : out  STD_LOGIC_VECTOR (0 to 10));
end prom_DMH;

architecture prom_DMH of prom_DMH is


constant ADDR_WIDTH: integer:=9;
constant DATA_WIDTH: integer:=11;

signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);

type rom_array is array (0 to 447)
        of std_logic_vector(DATA_WIDTH-1 downto 0);

constant rom: rom_array := (
	--x00 - cijfer_0
	"00111111100",    --0
	"01000000010",    --1
	"10000000001",    --2
	"10000000001",    --3
	"10000000001",    --4
	"10000000001",    --5
	"10000000001",    --6
	"10000000001",    --7
	"10000000001",    --8
	"10000000001",    --9
	"10000000001",    --10
	"10000000001",    --11
	"10000000001",    --12
	"10000000001",    --13
	"01000000010",    --14
	"00111111100",    --15
	
	
	--x01 - cijfer_1
	"00000000001",    --1
	"00000000001",    --1
	"00000000001",    --2
	"00000000001",    --3
	"00000000001",    --4
	"00000000001",    --5
	"00000000001",    --6
	"00000000001",    --7
	"00000000001",    --8
	"00000000001",    --9
	"00000000001",    --10
	"00000000001",    --11
	"00000000001",    --12
	"00000000001",    --13
	"00000000001",    --14
	"00000000001",    --15
	
	--x02 - cijfer_2
	"01111111100",    --1
	"00000000010",    --1
	"00000000001",    --2
	"00000000001",    --3
	"00000000001",    --4
	"00000000001",    --5
	"00000000010",    --6
	"00111111100",    --7
	"01000000000",    --8
	"10000000000",    --9
	"10000000000",    --10
	"10000000000",    --11
	"10000000000",    --12
	"10000000000",    --13
	"01000000000",    --14
	"00111111110",    --15
	
	--x03 - cijfer_3
	"11111111100",    --1
	"00000000010",    --1
	"00000000001",    --2
	"00000000001",    --3
	"00000000001",    --4
	"00000000001",    --5
	"00000000001",    --6
	"11111111111",    --7
	"00000000001",    --8
	"00000000001",    --9
	"00000000001",    --10
	"00000000001",    --11
	"00000000001",    --12
	"00000000001",    --13
	"00000000010",    --14
	"11111111100",    --15
	
	--x04 - cijfer_4
	"10000000001",	  --0
	"10000000001",    --1
	"10000000001",    --2
	"10000000001",    --3
	"10000000001",    --4
	"10000000001",    --5
	"01000000011",    --6
	"00111111101",    --7
	"00000000001",    --8
	"00000000001",    --9
	"00000000001",    --10
	"00000000001",    --11
	"00000000001",    --12
	"00000000001",    --13
	"00000000001",    --14
	"00000000001",    --15
	
	--x05 - cijfer_5
	"00111111110",	  --0
	"01000000000",    --1
	"10000000000",    --2
	"10000000000",    --3
	"10000000000",    --4
	"10000000000",    --5
	"01000000000",    --6
	"00111111100",    --7
	"00000000010",    --8
	"00000000001",    --9
	"00000000001",    --10
	"00000000001",    --11
	"00000000001",    --12
	"00000000001",    --13
	"00000000010",    --14
	"01111111100",    --15
	
	--x06 - cijfer_6
	"00111111110",    --0
	"01000000000",	  --1
	"10000000000",    --2
	"10000000000",    --3
	"10000000000",    --4
	"10000000000",    --5
	"10000000000",    --6
	"10111111100",    --7
	"11000000010",    --8
	"10000000001",    --9
	"10000000001",    --10
	"10000000001",    --11
	"10000000001",    --12
	"10000000001",    --13
	"01000000010",    --14
	"00111111100",    --15
	
	--x07 - cijfer_7
	"11111111100",    --0
	"00000000010",    --1
	"00000000001",    --2
	"00000000001",    --3
	"00000000001",    --4
	"00000000001",    --5
	"00000000001",    --6
	"00000000001",    --7
	"00000000001",    --8
	"00000000001",    --9
	"00000000001",    --10
	"00000000001",    --11
	"00000000001",    --12
	"00000000001",    --13
	"00000000001",    --14
	"00000000001",    --15
	
	--x08 - cijfer_8
	"00111111100",    --0
	"01000000010",	  --1
	"10000000001",    --2
	"10000000001",    --3
	"10000000001",    --4
	"10000000001",    --5
	"10000000001",    --6
	"11111111111",    --7
	"10000000001",    --8
	"10000000001",    --9
	"10000000001",    --10
	"10000000001",    --11
	"10000000001",    --12
	"10000000001",    --13
	"01000000010",    --14
	"00111111100",    --15
	
	--x09 - cijfer_9
	"00111111100",    --0
	"01000000010",    --1
	"10000000001",    --2
	"10000000001",    --3
	"10000000001",    --4
	"10000000001",    --5
	"01000000011",    --6
	"00111111101",    --7
	"00000000001",    --8
	"00000000001",    --9
	"00000000001",    --10
	"00000000001",    --11
	"00000000001",    --12
	"00000000001",    --13
	"00000000010",    --14
	"01111111100",    --15
	
	--x0a - zero
	"00000000000",    --0
	"00000000000",    --1
	"00000000000",    --2
	"00000000000",    --3
	"00000000000",    --4
	"00000000000",    --5
	"00000000000",    --6
	"00000000000",    --7
	"00000000000",    --8
	"00000000000",    --9
	"00000000000",    --10
	"00000000000",    --11
	"00000000000",    --12
	"00000000000",    --13
	"00000000000",    --14
	"00000000000",    --15
	
	--x0b - letter_a
	"11111111111",	 --0
	"10000000001",    --1
	"10000000001",    --2
	"10000000001",    --3
	"10000000001",    --4
	"10000000001",    --5
	"11111111111",    --6
	"10000000001",    --7
	"10000000001",    --8
	"10000000001",    --9
	"10000000001",    --10
	"10000000001",    --11
	"10000000001",    --12
	"10000000001",    --13
	"10000000001",    --14
	"10000000001",    --15
	
	--x0c - letter_c
	"11111111111",	 --0
	"10000000000",    --1
	"10000000000",    --2
	"10000000000",    --3
	"10000000000",    --4
	"10000000000",    --5
	"10000000000",    --6
	"10000000000",    --7
	"10000000000",    --8
	"10000000000",    --9
	"10000000000",    --10
	"10000000000",    --11
	"10000000000",    --12
	"10000000000",    --13
	"10000000000",    --14
	"11111111111",    --15
	
	--x0d - letter d
	"11111110000",	 --0
	"10000001000",    --1
	"10000000100",    --2
	"10000000010",    --3
	"10000000001",    --4
	"10000000001",    --5
	"10000000001",    --6
	"10000000001",    --7
	"10000000001",    --8
	"10000000001",    --9
	"10000000001",    --10
	"10000000001",    --11
	"10000000010",    --12
	"10000000100",    --13
	"10000001000",    --14
	"11111110000",    --15
	
	--x0e - letter e
	"11111111111",	 --0
	"10000000000", 	 --1
	"10000000000",    --2
	"10000000000",    --3
	"10000000000",    --4
	"10000000000",    --5
	"10000000000",    --6
	"11111111111",    --7
	"10000000000",    --8
	"10000000000",    --9
	"10000000000",    --10
	"10000000000",    --11
	"10000000000",    --12
	"10000000000",    --13
	"10000000000",    --14
	"11111111111",    --15
	
	--x0f - letter_h
	"10000000001",    --0
	"10000000001",    --1
	"10000000001",    --2
	"10000000001",    --3
	"10000000001",    --4
	"10000000001",    --5
	"10000000001",    --6
	"11111111111",    --7
	"10000000001",    --8
	"10000000001",    --9
	"10000000001",    --10
	"10000000001",    --11
	"10000000001",    --12
	"10000000001",    --13
	"10000000001",    --14
	"10000000001",    --15
	
	--x10 - letter_i
	"00000100000",    --0
	"00000100000",    --1
	"00000000000",    --2
	"00000100000",    --3
	"00000100000",    --4
	"00000100000",    --5
	"00000100000",    --6
	"00000100000",    --7
	"00000100000",    --8
	"00000100000",    --9
	"00000100000",    --10
	"00000100000",    --11
	"00000100000",    --12
	"00000100000",    --13
	"00000100000",    --14
	"00000100000",    --15
	
	--x11 - letter_j
	"00000100000",    --0
	"00000100000",    --1
	"00000000000",    --2
	"00000100000",    --3
	"00000100000",    --4
	"00000100000",    --5
	"00000100000",    --6
	"00000100000",    --7
	"00000100000",    --8
	"00000100000",    --9
	"00000100000",    --10
	"00000100000",    --11
	"10000100000",    --12
	"10000100000",    --13
	"01001000000",    --14
	"00110000000",    --15
	
	--x12 - letter_k
	"10000000001",    --0
	"10000000010",    --1
	"10000000100",    --2
	"10000001000",    --3
	"10000010000",    --4
	"10000100000",    --5
	"10001000000",    --6
	"11110000000",    --7
	"11110000000",    --8
	"10001000000",    --9
	"10000100000",    --10
	"10000010000",    --11
	"10000001000",    --12
	"10000000100",    --13
	"10000000010",    --14
	"10000000001",    --15
	
	--x13 - letter_m
	"10000000001",    --0
	"11000000011",    --1
	"10100000101",    --2
	"10010001001",    --3
	"10001010001",    --4
	"10000100001",    --5
	"10000000001",    --6
	"10000000001",    --7
	"10000000001",    --8
	"10000000001",    --9
	"10000000001",    --10
	"10000000001",    --11
	"10000000001",    --12
	"10000000001",    --13
	"10000000001",    --14
	"10000000001",    --15
	
	--x14 - letter_n
	"10000000001",    --0
	"10000000001",    --1
	"10000000001",    --2
	"11000000001",    --3
	"10100000001",    --4
	"10010000001",    --5
	"10001000001",    --6
	"10000100001",    --7
	"10000010001",    --8
	"10000001001",    --9
	"10000000101",    --10
	"10000000011",    --11
	"10000000001",    --12
	"10000000001",    --13
	"10000000001",    --14
	"10000000001",    --15
	
	--x15 - letter_o
	"00111111100",    --0
	"01000000010",    --1
	"10000000001",    --2
	"10000000001",    --3
	"10000000001",    --4
	"10000000001",    --5
	"10000000001",    --6
	"10000000001",    --7
	"10000000001",    --8
	"10000000001",    --9
	"10000000001",    --10
	"10000000001",    --11
	"10000000001",    --12
	"10000000001",    --13
	"01000000010",    --14
	"00111111100",    --15
	
	--x16 - letter_r
	"11111111100",    --0
	"10000000010",    --1
	"10000000001",    --2
	"10000000001",    --3
	"10000000001",    --4
	"10000000001",    --5
	"10000000010",    --6
	"11111111100",    --7
	"10010000000",    --8
	"10001000000",    --9
	"10000100000",    --10
	"10000010000",    --11
	"10000001000",    --12
	"10000000100",    --13
	"10000000010",    --14
	"10000000001",    --15
	
	--x17 - letter_t
	"11111111111",    --0
	"00000100000",    --1
	"00000100000",    --2
	"00000100000",    --3
	"00000100000",    --4
	"00000100000",    --5
	"00000100000",    --6
	"00000100000",    --7
	"00000100000",    --8
	"00000100000",    --9
	"00000100000",    --10
	"00000100000",    --11
	"00000100000",    --12
	"00000100000",    --13
	"00000100000",    --14
	"00000100000",    --15
	
	--x18 - letter_u
	"10000000001",    --0
	"10000000001",    --1
	"10000000001",    --2
	"10000000001",    --3
	"10000000001",    --4
	"10000000001",    --5
	"10000000001",    --6
	"10000000001",    --7
	"10000000001",    --8
	"10000000001",    --9
	"10000000001",    --10
	"10000000001",    --11
	"10000000001",    --12
	"10000000001",    --13
	"10000000001",    --14
	"11111111111",    --15
	
	--x19 - letter_w
	"10000000001",    --0
	"10000000001",    --1
	"10000000001",    --2
	"10000000001",    --3
	"10000000001",    --4
	"10000000001",    --5
	"10000000001",    --6
	"10000000001",    --7
	"10000100001",    --8
	"10001010001",    --9
	"10010001001",    --10
	"10010001001",    --11
	"10100000101",    --12
	"10100000101",    --13
	"11000000011",    --14
	"10000000001",    --15
	
	--x1a - dubbele_punt
	"00000000000",    --0
	"00000000000",    --1
	"00000000000",    --2
	"00001110000",    --3
	"00001110000",    --4
	"00001110000",    --5
	"00000000000",    --6
	"00000000000",    --7
	"00000000000",    --8
	"00000000000",    --9
	"00001110000",    --10
	"00001110000",    --11
	"00001110000",    --12
	"00000000000",    --13
	"00000000000",   --14
	"00000000000",    --15
	
	
	--x1b - schuine_streep
	"00000000001",    --0
	"00000000011",    --1
	"00000000010",    --2
	"00000000100",    --3
	"00000000100",    --4
	"00000001000",    --5
	"00000001000",    --6
	"00000010000",    --7
	"00000010000",    --8
	"00000100000",    --9
	"00000100000",    --10
	"00001000000",    --11
	"00001000000",    --12
	"00010000000",    --13
	"00010000000",    --14
	"00100000000"     --15
	
);

begin

	process (clk)
   begin
      if rising_edge(clk) then
        addr_reg <= addr;
      end if;
   end process;
	M <= ROM(conv_integer(unsigned(addr_reg)));
	
end prom_DMH;

