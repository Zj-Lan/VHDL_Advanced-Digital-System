LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY fpq IS
	PORT(clk:IN STD_LOGIC;
	clk_out:OUT STD_LOGIC);
END fpq;

ARCHITECTURE dwz OF fpq IS

	CONSTANT m : INTEGER:=2;
	SIGNAL tmp :STD_LOGIC;

	BEGIN

	PROCESS(clk, tmp)
	VARIABLE cout : INTEGER:=0;
	
	BEGIN
		IF clk'EVENT AND clk='1' THEN cout:=cout+1;
			IF cout<=m THEN tmp<='0';
			ELSIF cout<m*2 THEN tmp<='1';
			ELSE cout:=0;	
			END IF;
		END IF;
		
	END PROCESS;
	clk_out<=tmp;
END dwz;